// Reference from week6 lab2 module.
package bus_trans_pkg;
    typedef enum  {READ, WRITE} op_kind_e;
    `include "bus_trans.sv"
    `include "drived_trans.sv"

endpackage